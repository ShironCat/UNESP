-- megafunction wizard: %RAM: 1-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: RAM1Port.vhd
-- Megafunction Name(s):
-- 			altsyncram
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 350 03/24/2010 SP 2 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY RAM1Port IS
	PORT
	(
		iSW		 : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
		iKEY	 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
		q		 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		oHEX0_D  : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		oHEX0_DP : OUT STD_LOGIC;
		oHEX1_D  : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		oHEX1_DP : OUT STD_LOGIC;
		oHEX2_D  : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		oHEX2_DP : OUT STD_LOGIC
	);
END RAM1Port;


ARCHITECTURE SYN OF ram1port IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	--SIGNAL q			: STD_LOGIC_VECTOR (3 DOWNTO 0);


	COMPONENT altsyncram
	GENERIC (
		clock_enable_input_a		: STRING;
		clock_enable_output_a		: STRING;
		intended_device_family		: STRING;
		lpm_hint		            : STRING;
		lpm_type		            : STRING;
		numwords_a		            : NATURAL;
		operation_mode				: STRING;
		outdata_aclr_a				: STRING;
		outdata_reg_a				: STRING;
		power_up_uninitialized		: STRING;
		ram_block_type				: STRING;
		widthad_a					: NATURAL;
		width_a						: NATURAL;
		width_byteena_a				: NATURAL
	);
	PORT (
			wren_a		: IN STD_LOGIC_VECTOR( 0 downto 0);
			clock0		: IN STD_LOGIC_VECTOR( 0 downto 0);
			address_a	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			q_a			: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			data_a		: IN STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
	END COMPONENT;

	COMPONENT BinToHex4 is
	PORT (
	iSW      : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	oHEX0_D  : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	oHEX0_DP : OUT STD_LOGIC
	);
	END COMPONENT;

BEGIN
	q    <= sub_wire0(3 DOWNTO 0);

	altsyncram_component : altsyncram
	GENERIC MAP (
		clock_enable_input_a => "BYPASS",
		clock_enable_output_a => "BYPASS",
		intended_device_family => "Cyclone II",
		lpm_hint => "ENABLE_RUNTIME_MOD=NO",
		lpm_type => "altsyncram",
		numwords_a => 16,
		operation_mode => "SINGLE_PORT",
		outdata_aclr_a => "NONE",
		outdata_reg_a => "UNREGISTERED",
		power_up_uninitialized => "FALSE",
		ram_block_type => "M4K",
		widthad_a => 4,
		width_a => 4,
		width_byteena_a => 1
	)
	PORT MAP (
		wren_a => iSW(8 DOWNTO 8),
		clock0 => iKEY(0 DOWNTO 0),
		address_a => iSW(3 DOWNTO 0),
		data_a => iSW(7 DOWNTO 4),
		q_a => sub_wire0
	);

	--Endere�o
	bin1: BinToHex4 port map(iSW(3 DOWNTO 0), oHEX0_D(6 DOWNTO 0), oHEX0_DP);
	--Dados de entrada
	bin2: BinToHex4 port map(iSW(7 DOWNTO 4), oHEX1_D(6 DOWNTO 0), oHEX1_DP);
	--Dados de sa�da
	bin3: BinToHex4 port map(sub_wire0(3 DOWNTO 0), oHEX2_D(6 DOWNTO 0), oHEX2_DP);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADDRESSSTALL_A NUMERIC "0"
-- Retrieval info: PRIVATE: AclrAddr NUMERIC "0"
-- Retrieval info: PRIVATE: AclrByte NUMERIC "0"
-- Retrieval info: PRIVATE: AclrData NUMERIC "0"
-- Retrieval info: PRIVATE: AclrOutput NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_ENABLE NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_SIZE NUMERIC "8"
-- Retrieval info: PRIVATE: BlankMemory NUMERIC "1"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_A NUMERIC "0"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_A NUMERIC "0"
-- Retrieval info: PRIVATE: Clken NUMERIC "0"
-- Retrieval info: PRIVATE: DataBusSeparated NUMERIC "1"
-- Retrieval info: PRIVATE: IMPLEMENT_IN_LES NUMERIC "0"
-- Retrieval info: PRIVATE: INIT_FILE_LAYOUT STRING "PORT_A"
-- Retrieval info: PRIVATE: INIT_TO_SIM_X NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: PRIVATE: JTAG_ENABLED NUMERIC "0"
-- Retrieval info: PRIVATE: JTAG_ID STRING "NONE"
-- Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
-- Retrieval info: PRIVATE: MIFfilename STRING ""
-- Retrieval info: PRIVATE: NUMWORDS_A NUMERIC "16"
-- Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "2"
-- Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_A NUMERIC "3"
-- Retrieval info: PRIVATE: RegAddr NUMERIC "1"
-- Retrieval info: PRIVATE: RegData NUMERIC "1"
-- Retrieval info: PRIVATE: RegOutput NUMERIC "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: SingleClock NUMERIC "1"
-- Retrieval info: PRIVATE: UseDQRAM NUMERIC "1"
-- Retrieval info: PRIVATE: WRCONTROL_ACLR_A NUMERIC "0"
-- Retrieval info: PRIVATE: WidthAddr NUMERIC "4"
-- Retrieval info: PRIVATE: WidthData NUMERIC "4"
-- Retrieval info: PRIVATE: rden NUMERIC "0"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_A STRING "BYPASS"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_A STRING "BYPASS"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: CONSTANT: LPM_HINT STRING "ENABLE_RUNTIME_MOD=NO"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altsyncram"
-- Retrieval info: CONSTANT: NUMWORDS_A NUMERIC "16"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "SINGLE_PORT"
-- Retrieval info: CONSTANT: OUTDATA_ACLR_A STRING "NONE"
-- Retrieval info: CONSTANT: OUTDATA_REG_A STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: POWER_UP_UNINITIALIZED STRING "FALSE"
-- Retrieval info: CONSTANT: RAM_BLOCK_TYPE STRING "M4K"
-- Retrieval info: CONSTANT: WIDTHAD_A NUMERIC "4"
-- Retrieval info: CONSTANT: WIDTH_A NUMERIC "4"
-- Retrieval info: CONSTANT: WIDTH_BYTEENA_A NUMERIC "1"
-- Retrieval info: USED_PORT: address 0 0 4 0 INPUT NODEFVAL address[3..0]
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT VCC clock
-- Retrieval info: USED_PORT: data 0 0 4 0 INPUT NODEFVAL data[3..0]
-- Retrieval info: USED_PORT: q 0 0 4 0 OUTPUT NODEFVAL q[3..0]
-- Retrieval info: USED_PORT: wren 0 0 0 0 INPUT NODEFVAL wren
-- Retrieval info: CONNECT: @address_a 0 0 4 0 address 0 0 4 0
-- Retrieval info: CONNECT: q 0 0 4 0 @q_a 0 0 4 0
-- Retrieval info: CONNECT: @clock0 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @data_a 0 0 4 0 data 0 0 4 0
-- Retrieval info: CONNECT: @wren_a 0 0 0 0 wren 0 0 0 0
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL RAM1Port.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL RAM1Port.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL RAM1Port.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL RAM1Port.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL RAM1Port_inst.vhd FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL RAM1Port_waveforms.html TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL RAM1Port_wave*.jpg FALSE
-- Retrieval info: LIB_FILE: altera_mf
