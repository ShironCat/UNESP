LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY BinToHex8 IS
PORT (
	iSW : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	oHEX0_D : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	oHEX1_D : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
	oHEX0_DP : OUT STD_LOGIC;
	oHEX1_DP : OUT STD_LOGIC
);
END BinToHex8;

ARCHITECTURE BinToHex8Comportamento OF BinToHex8 IS
COMPONENT BinToHex4 is 
	PORT (
	iSW : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	oHEX0_D : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	oHEX0_DP : OUT STD_LOGIC
);
END COMPONENT;
BEGIN
	display1 : BinToHex4 port map(iSW(3 DOWNTO 0), oHEX0_D, oHEX0_DP);
	display2 : BinToHex4 port map(iSW(7 DOWNTO 4), oHEX1_D, oHEX1_DP);
END BinToHex8Comportamento;